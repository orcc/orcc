-------------------------------------------------------------------------------
-- Title      : BroadCast
-- Project    : ORCC
-------------------------------------------------------------------------------
-- File       : broadcast.vhd
-- Author     : Nicolas Siret (nicolas.siret@live.fr)
-- Company    : Lead Tech Design
-- Created    : 
-- Last update: 2011-02-02
-- Platform   : 
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Copyright (c) 2009-2010, LEAD TECH DESIGN Rennes - France
-- Copyright (c) 2009-2010, IETR/INSA of Rennes
-- All rights reserved.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--  -- Redistributions of source code must retain the above copyright notice,
--     this list of conditions and the following disclaimer.
--  -- Redistributions in binary form must reproduce the above copyright notice,
--     this list of conditions and the following disclaimer in the documentation
--     and/or other materials provided with the distribution.
--  -- Neither the name of the IETR/INSA of Rennes nor the names of its
--     contributors may be used to endorse or promote products derived from this
--     software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY
-- WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2010-02-09  1.0      Nicolas      Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity broadcast is
  generic
    (
      width : integer := 16;
      size  : integer := 2);
  port
    (
      reset_n     : in  std_logic;
      clock       : in  std_logic;
      --
      input_data  : in  std_logic_vector (width -1 downto 0);
      input_send  : in  std_logic;
      input_ack   : out std_logic;
      --
      output_data : out std_logic_vector (width -1 downto 0);
      output_send : out std_logic_vector (size -1 downto 0);
      output_ack  : in  std_logic_vector (size -1 downto 0)
      );
end broadcast;


-------------------------------------------------------------------------------


architecture arch_broadcast of broadcast is

-------------------------------------------------------------------------------
-- Signals and constants declaration
-----------------------------------------------------------------------------
  constant ones        : std_logic_vector (size -1 downto 0) := (others => '1');
  --
  signal   internalAck : std_logic_vector (size -1 downto 0);
  
begin

  output_data <= input_data;

  -- Management of the external SEND (destination actor)
  externalSend : for i in 0 to size -1 generate
    output_send(i) <= input_send and not internalAck(i);
  end generate externalSend;


  -- Management of the external ACK (source actor)
  externalAck : process (output_ack, internalAck, input_send) is
  begin
    if ((output_ack or internalAck) = ones) then
      input_ack <= '1';
    else
      input_ack <= '0';
    end if;
  end process externalAck;

  
  -- Management of the internal ACK (source actor)
  counterGen : for i in 0 to size -1 generate
    process (clock, reset_n) is
    begin
      if reset_n = '0' then
        internalAck(i) <= '0';
      elsif rising_edge (clock) then
        if ((output_ack or internalAck) = ones) then
          internalAck(i) <= '0';
        elsif output_ack(i) = '1' then
          internalAck(i) <= '1';
        end if;
      end if;
    end process;
  end generate counterGen;
  
end arch_broadcast;

--------------------------------------------------------------------------
